use work.cfuncs.all;

entity tb is
end tb;

architecture arch of tb is
begin
  process begin
    hello_world;
    wait;
  end process;
end;
